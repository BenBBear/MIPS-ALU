library verilog;
use verilog.vl_types.all;
entity TESTmux_5bit is
end TESTmux_5bit;
