library verilog;
use verilog.vl_types.all;
entity TESTnot_32bit is
end TESTnot_32bit;
