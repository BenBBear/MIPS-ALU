module bitSlice_1bit (Out, Cout, A, B,Cin,Cntrl)
  input A,B,Cin;
  input [2:0] Cntrl;
  output Out, Cout;
  
endmodule
