library verilog;
use verilog.vl_types.all;
entity TESTadd_1bit is
end TESTadd_1bit;
