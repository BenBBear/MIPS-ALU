library verilog;
use verilog.vl_types.all;
entity TESTbitSlice_1bit is
end TESTbitSlice_1bit;
