`define NOT not #10

module not_32bit(in0,in1,in2,in3,in4,in5,in6,in7,in8,in9,in10,in11,in12,in13,in14,in15,in16,
                  in17,in18,in19,in20,in21,in22,in23,in24,in25,in26,in27,in28,in29,in30,in31,
                  out0,out1,out2,out3,out4,out5,out6,out7,out8,out9,out10,out11,out12,out13,
                  out14,out15,out16,out17,out18,out19,out20,out21,out22,out23,out24,out25,
                  out26,out27,out28,out29,out30,out31);
  input in0,in1,in2,in3,in4,in5,in6,in7,in8,in9,in10,in11,in12,in13,in14,in15,in16,
          in17,in18,in19,in20,in21,in22,in23,in24,in25,in26,in27,in28,in29,in30,in31;
  output out0,out1,out2,out3,out4,out5,out6,out7,out8,out9,out10,out11,out12,out13,
          out14,out15,out16,out17,out18,out19,out20,out21,out22,out23,out24,out25,
          out26,out27,out28,out29,out30,out31;

  `NOT not0(out0,in0);
  `NOT not1(out1,in1);
  `NOT not2(out2,in2);
  `NOT not3(out3,in3);
  `NOT not4(out4,in4);
  `NOT not5(out5,in5);
  `NOT not6(out6,in6);
  `NOT not7(out7,in7);
  `NOT not8(out8,in8);
  `NOT not9(out9,in9);
  `NOT not10(out10,in10);
  `NOT not11(out11,in11);
  `NOT not12(out12,in12);
  `NOT not13(out13,in13);
  `NOT not14(out14,in14);
  `NOT not15(out15,in15);
  `NOT not16(out16,in16);
  `NOT not17(out17,in17);
  `NOT not18(out18,in18);
  `NOT not19(out19,in19);
  `NOT not20(out20,in20);
  `NOT not21(out21,in21);
  `NOT not22(out22,in22);
  `NOT not23(out23,in23);
  `NOT not24(out24,in24);
  `NOT not25(out25,in25);
  `NOT not26(out26,in26);
  `NOT not27(out27,in27);
  `NOT not28(out28,in28);
  `NOT not29(out29,in29);
  `NOT not30(out30,in30);
  `NOT not31(out31,in31);
endmodule